package Tb;

import MMTED::*;
import StmtFSM::*;
import Complex::*;
import FixedPoint::*;

(* synthesize *)
module mkTb (Empty);
    MMTED_IFC mmTed <- mkMMTED;
 
    Stmt test = seq
        mmTed.addSample(cmplx(0.00000045 , 0.00000000));
        mmTed.addSample(cmplx(-0.00000063 , -0.00000000));
        mmTed.addSample(cmplx(0.00000176 , 0.00000000));
        mmTed.addSample(cmplx(-0.00000105 , -0.00000000));
        mmTed.addSample(cmplx(0.00000404 , 0.00000000));
        mmTed.addSample(cmplx(-0.00000582 , -0.00000000));
        mmTed.addSample(cmplx(0.00000486 , 0.00000000));
        mmTed.addSample(cmplx(-0.00001356 , -0.00000000));
        mmTed.addSample(cmplx(0.00001463 , 0.00000000));
        mmTed.addSample(cmplx(-0.00002411 , -0.00000000));
        mmTed.addSample(cmplx(0.00005032 , 0.00000000));
        mmTed.addSample(cmplx(-0.00060910 , -0.00000000));
        mmTed.addSample(cmplx(-0.00006652 , -0.00000000));
        mmTed.addSample(cmplx(-0.00063801 , -0.00000000));
        mmTed.addSample(cmplx(-0.00247127 , -0.00000000));
        mmTed.addSample(cmplx(-0.00231275 , -0.00000000));
        mmTed.addSample(cmplx(-0.00030051 , -0.00000000));
        mmTed.addSample(cmplx(0.00447211 , 0.00000000));
        mmTed.addSample(cmplx(0.00813003 , 0.00000000));
        mmTed.addSample(cmplx(0.00519995 , 0.00000000));
        mmTed.addSample(cmplx(0.00004130 , 0.00000000));
        mmTed.addSample(cmplx(-0.00104713 , -0.00000000));
        mmTed.addSample(cmplx(0.00758543 , 0.00000000));
        mmTed.addSample(cmplx(0.01650484 , 0.00000000));
        mmTed.addSample(cmplx(0.00382114 , 0.00000000));
        mmTed.addSample(cmplx(-0.05110755 , -0.00000000));
        mmTed.addSample(cmplx(-0.12753011 , -0.00000000));
        mmTed.addSample(cmplx(-0.15057974 , -0.00000000));
        mmTed.addSample(cmplx(-0.02356299 , -0.00000000));
        mmTed.addSample(cmplx(0.28862881 , 0.00000000));
        mmTed.addSample(cmplx(0.70031729 , 0.00000000));
        mmTed.addSample(cmplx(1.01521421 , 0.00000000));
        mmTed.addSample(cmplx(1.02095187 , 0.00000000));
        mmTed.addSample(cmplx(0.63395561 , 0.00000000));
        mmTed.addSample(cmplx(-0.02441158 , -0.00000000));
        mmTed.addSample(cmplx(-0.66884167 , -0.00000000));
        mmTed.addSample(cmplx(-0.99340829 , -0.00000000));
        mmTed.addSample(cmplx(-0.84519362 , -0.00000000));
        mmTed.addSample(cmplx(-0.29898719 , -0.00000000));
        mmTed.addSample(cmplx(0.39654926 , 0.00000000));
        mmTed.addSample(cmplx(0.95945283 , 0.00000000));
        mmTed.addSample(cmplx(1.22849398 , 0.00000000));
        mmTed.addSample(cmplx(1.21996377 , 0.00000000));
        mmTed.addSample(cmplx(1.08610143 , 0.00000000));
        mmTed.addSample(cmplx(1.00061948 , 0.00000000));
        mmTed.addSample(cmplx(1.05329518 , 0.00000000));
        mmTed.addSample(cmplx(1.19003194 , 0.00000000));
        mmTed.addSample(cmplx(1.24266932 , 0.00000000));
        mmTed.addSample(cmplx(1.03865105 , 0.00000000));
        mmTed.addSample(cmplx(0.51862961 , 0.00000000));
        mmTed.addSample(cmplx(-0.18542223 , -0.00000000));
        mmTed.addSample(cmplx(-0.78956960 , -0.00000000));
        mmTed.addSample(cmplx(-1.00554118 , -0.00000000));
        mmTed.addSample(cmplx(-0.71469196 , -0.00000000));
        mmTed.addSample(cmplx(-0.05891549 , -0.00000000));
        mmTed.addSample(cmplx(0.62431948 , 0.00000000));
        mmTed.addSample(cmplx(0.98971031 , 0.00000000));
        mmTed.addSample(cmplx(0.86987467 , 0.00000000));
        mmTed.addSample(cmplx(0.34365957 , 0.00000000));
        mmTed.addSample(cmplx(-0.34615171 , -0.00000000));
        mmTed.addSample(cmplx(-0.95104756 , -0.00000000));
        mmTed.addSample(cmplx(-1.32933262 , -0.00000000));
        mmTed.addSample(cmplx(-1.45512862 , -0.00000000));
        mmTed.addSample(cmplx(-1.35307716 , -0.00000000));
        mmTed.addSample(cmplx(-1.04180801 , -0.00000000));
        mmTed.addSample(cmplx(-0.54267257 , -0.00000000));
        mmTed.addSample(cmplx(0.06757424 , 0.00000000));
        mmTed.addSample(cmplx(0.63496489 , 0.00000000));
        mmTed.addSample(cmplx(0.98227945 , 0.00000000));
        mmTed.addSample(cmplx(1.00723280 , 0.00000000));
        mmTed.addSample(cmplx(0.74708594 , 0.00000000));
        mmTed.addSample(cmplx(0.35827650 , 0.00000000));
        mmTed.addSample(cmplx(0.02450761 , 0.00000000));
        mmTed.addSample(cmplx(-0.14432827 , -0.00000000));
        mmTed.addSample(cmplx(-0.15123293 , -0.00000000));
        mmTed.addSample(cmplx(-0.07592963 , -0.00000000));
        mmTed.addSample(cmplx(-0.00464254 , -0.00000000));
        mmTed.addSample(cmplx(0.02283014 , 0.00000000));
        mmTed.addSample(cmplx(0.01597087 , 0.00000000));
        mmTed.addSample(cmplx(0.00258442 , 0.00000000));
        mmTed.addSample(cmplx(-0.00014104 , -0.00000000));
        mmTed.addSample(cmplx(0.00512518 , 0.00000000));
        mmTed.addSample(cmplx(0.00828380 , 0.00000000));
        mmTed.addSample(cmplx(0.00550764 , 0.00000000));
        mmTed.addSample(cmplx(0.00040432 , 0.00000000));
        mmTed.addSample(cmplx(-0.00273708 , -0.00000000));
        mmTed.addSample(cmplx(-0.00272784 , -0.00000000));
        mmTed.addSample(cmplx(-0.00099175 , -0.00000000));
        mmTed.addSample(cmplx(-0.00002388 , -0.00000000));
        mmTed.addSample(cmplx(0.00000417 , 0.00000000));
        mmTed.addSample(cmplx(-0.00000044 , -0.00000000));
        mmTed.addSample(cmplx(0.00000458 , 0.00000000));
        mmTed.addSample(cmplx(0.00000267 , 0.00000000));
        mmTed.addSample(cmplx(0.00000126 , 0.00000000));
        mmTed.addSample(cmplx(-0.00000127 , -0.00000000));
        mmTed.addSample(cmplx(-0.00000126 , -0.00000000));
        mmTed.addSample(cmplx(-0.00000076 , -0.00000000));
        mmTed.addSample(cmplx(-0.00000000 , -0.00000000));
        mmTed.addSample(cmplx(0.00000000 , 0.00000000));
        mmTed.addSample(cmplx(0.00000000 , 0.00000000));
        mmTed.addSample(cmplx(0.00000000 , 0.00000000));
        $write("timing error: ");
        action
        let err <- mmTed.getError;
        fxptWrite(5,err);
        endaction
        $display("  ");
    endseq;
    mkAutoFSM(test);
    
endmodule: mkTb
endpackage: Tb
