package FIRcoeff;

typedef Int#(13) Sample_Type;
Integer n_TAPS = 43;

Sample_Type coeff[n_TAPS] ={186, 233, 248, 217, 134, 0, -173, -364, -540, -665, 
-700, -613, -382, 0, 521, 1151, 1842, 2533, 3159, 3660, 3983, 4095, 3983, 3660,
3159, 2533, 1842, 1151, 521, 0, -382, -613, -700, -665, -540, -364, -173, 0,  
134,  217,  248,  233, 186};

endpackage: FIRcoeff
