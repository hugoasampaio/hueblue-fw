package FIRcoeff;
import FixedPoint::*;

//typedef FixedPoint#(3, 32) FIRtap_Type;
//typedef Real FIRtap_Type;
typedef Int#(16) FIRtap_Type;
Integer n_TAPS = 43;


FIRtap_Type coeff[n_TAPS] ={186, 233, 248, 217, 134, 0, -173, -364, -540, -665, 
-700, -613, -382, 0, 521, 1151, 1842, 2533, 3159, 3660, 3983, 4095, 3983, 3660,
3159, 2533, 1842, 1151, 521, 0, -382, -613, -700, -665, -540, -364, -173, 0,  
134,  217,  248,  233, 186};

/*
FIRtap_Type coeff[n_TAPS] = {
 -0.01897049, 
 -0.01842133, 
 -0.00954316,  
  0.00624239,  
  0.02459163,  
  0.03898283,
  0.04231734,  
  0.02906669, 
 -0.00255221, 
 -0.04897974, 
 -0.10083352, 
 -0.1438624,
 -0.16131922, 
 -0.13737078, 
 -0.0608575,   
  0.07144658,  
  0.25288767,  
  0.46687654,
  0.68890519,  
  0.89035557,  
  1.04339768,  
  1.12599805,  
  1.12599805,  
  1.04339768,
  0.89035557,  
  0.68890519,  
  0.46687654, 
  0.25288767,  
  0.07144658, 
 -0.0608575,
 -0.13737078, 
 -0.16131922, 
 -0.1438624,  
 -0.10083352, 
 -0.04897974, 
 -0.00255221,
  0.02906669,  
  0.04231734,  
  0.03898283,  
  0.02459163,  
  0.00624239, 
 -0.00954316,
 -0.01842133};
*/
endpackage: FIRcoeff
